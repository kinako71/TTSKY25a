VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TOP
  CLASS BLOCK ;
  FOREIGN TOP ;
  ORIGIN 0.855 1.275 ;
  SIZE 4.370 BY 5.070 ;
  OBS
      LAYER nwell ;
        RECT -0.855 1.525 3.515 3.395 ;
      LAYER pwell ;
        RECT -0.855 0.845 0.155 1.525 ;
      LAYER nwell ;
        RECT 0.155 0.845 3.515 1.525 ;
        RECT -0.855 -0.875 3.515 0.845 ;
      LAYER li1 ;
        RECT -0.660 -1.195 3.320 3.715 ;
      LAYER met1 ;
        RECT -0.720 -1.225 3.380 3.745 ;
  END
END TOP
END LIBRARY

